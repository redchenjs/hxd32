/*
 * core_config.sv
 *
 *  Created on: 2021-08-18 19:51
 *      Author: Jack Chen <redchenjs@live.com>
 */

`ifndef _CORE_CONFIG_SV_
`define _CORE_CONFIG_SV_

/* Base ISA */
`define CONFIG_ISA_RV32I

/* Extensions */
`define CONFIG_ISA_RV32C

`endif
